// -----------------------------------------------------------------------------
// zeropad_rows.v
//  - �Է�(mp) �� ������( W x HIN )�� ���� ĸó�ϸ鼭 mp_valid �޽� ������ ����
//  - �� ����(slot_period)�� TOP 4�� �� ĸó�� ��� 24�� �� BOT 4����
//    "mp_validó�� 1clk �޽�"�� ������ (���� ���� ���� ��ġ)
//  - ��� ����/������ ��赵 slot_period ������� ��Ȯ�� 1clk �޽�
//  - ���� �������� �ٽ� CAP �� TOP �� PAY �� BOT ��ȯ (1-������ �����Ͻ�)
// -----------------------------------------------------------------------------
`timescale 1ns/1ps
module zeropad_rows #(
  parameter integer W   = 32,
  parameter integer HIN = 24,
  parameter integer PAD = 4
)(
  input  wire       clk,
  input  wire       srst,            // active-HIGH

  // �Է�: mp �������� ��� (1�ȼ�/�޽�)
  input  wire       in_valid,        // mp_valid
  input  wire [7:0] in_pixel,        // mp_pixel
  input  wire       in_line_last,    // mp_line_last (�� �� ������ �ȼ����� 1clk)

  // ���: �е� ���� (W x (HIN+2*PAD))
  output reg        out_valid,
  output reg [7:0]  out_pixel,
  output reg        out_line_last,   // �� �� ������ �ȼ����� 1clk
  output reg        out_frame_last,  // ������ ������ �ȼ����� 1clk
  output reg        out_is_pad       // �е� ����(Top/Bot)���� 1
);

  // --------------------------
  // ��ƿ: ���� clog2 (Verilog-2001)
  // --------------------------
  function integer CLOG2;
    input integer x;
    integer i;
    begin
      i = 0;
      while ((1<<i) < x) i = i + 1;
      CLOG2 = i;
    end
  endfunction

  // --------------------------
  // ������ ���� (W*HIN ����Ʈ)
  // --------------------------
  localparam integer DEPTH = W*HIN;
  localparam integer A_W   = CLOG2(DEPTH);

  reg [7:0] fb [0:DEPTH-1];

  reg [A_W-1:0] wr_addr;      // CAP���� ���
  reg [A_W-1:0] rd_addr;      // PAY���� ���

  // --------------------------
  // ���� ���� (mp_valid �޽� ����)
  // --------------------------
  reg        iv_d;
  wire       iv_rise = in_valid & ~iv_d;

  reg        ill_d;
  wire       ill_rise = in_line_last & ~ill_d;

  reg [15:0] slot_cnt;
  reg [15:0] slot_period;     // ���� ���� �� mp_valid ����(Ŭ����)

  // --------------------------
  // ����/ī����
  // --------------------------
  localparam [2:0] S_CAP = 3'd0,  // �Է� ������ ĸó + ���� ����
                   S_TOP = 3'd1,  // TOP PAD  (PAD lines)
                   S_PAY = 3'd2,  // PAYLOAD  (HIN lines)
                   S_BOT = 3'd3;  // BOTTOM PAD (PAD lines)

  reg [2:0] st;

  // PAD/��� ���� ����(���� ����)
  reg [9:0] px_in_line;       // 0..W-1 (���� ���� ����)
  reg [6:0] lines_done;       // ������ ���� �� (Top/PAY/Bot �������� ���)

  // PAD/����� ���� ƽ (mp_valid ������ ������ ������ 1clk �޽�)
  reg  [15:0] gen_cnt;
  wire        have_tempo = (slot_period != 16'd0);
  wire        slot_tick  = have_tempo && (gen_cnt == slot_period - 1);

  // --------------------------
  // ���� ����
  // --------------------------
  integer i;
  always @(posedge clk) begin
    if (srst) begin
      // �Է��� edge �����
      iv_d        <= 1'b0;
      ill_d       <= 1'b0;

      // ���� ����
      slot_cnt    <= 16'd0;
      slot_period <= 16'd0;

      // ������ ���� �ּ�
      wr_addr     <= {A_W{1'b0}};
      rd_addr     <= {A_W{1'b0}};

      // ���/���� �ʱ�ȭ
      out_valid      <= 1'b0;
      out_pixel      <= 8'd0;
      out_line_last  <= 1'b0;
      out_frame_last <= 1'b0;
      out_is_pad     <= 1'b0;

      st          <= S_CAP;
      px_in_line  <= 10'd0;
      lines_done  <= 7'd0;
      gen_cnt     <= 16'd0;

    end else begin
      // edge ����� ����
      iv_d  <= in_valid;
      ill_d <= in_line_last;

      // �⺻ ��� ����Ʈ
      out_valid      <= 1'b0;
      out_line_last  <= 1'b0;
      out_frame_last <= 1'b0;
      out_is_pad     <= 1'b0;

      //------------------------------------------------------
      // ����(���� ����) ����: ���� ���� ������ in_valid ��� ������ ����
      //------------------------------------------------------
      slot_cnt <= slot_cnt + 16'd1;
      if (iv_rise) begin
        // ù �޽� �ĺ��� ���� ����
        if (slot_period == 16'd0)
          slot_period <= slot_cnt;     // �ʱⰪ
        else
          slot_period <= slot_cnt;     // �ʿ�� �̵���� ������ ����ȭ ����
        slot_cnt <= 16'd1;             // ���� �޽����� �ٽ� ���� ����
      end
      if (ill_rise) begin
        slot_cnt <= 16'd0;             // ���� �ѱ� �� ī���� �����
      end

      //------------------------------------------------------
      // PAD/����� ���� ƽ �߻���
      //------------------------------------------------------
      if (st==S_TOP || st==S_PAY || st==S_BOT) begin
        if (have_tempo) begin
          gen_cnt <= slot_tick ? 16'd0 : (gen_cnt + 16'd1);
        end else begin
          gen_cnt <= 16'd0; // ���� ��Ȯ���̸� ���
        end
      end else begin
        gen_cnt <= 16'd0;   // CAP������ ƽ ī���� ����
      end

      //------------------------------------------------------
      // ���±��
      //------------------------------------------------------
      case (st)
        // ====================================================
        // 1) CAPTURE (�Է� ������ ��ü ���� + ���� ����)
        // ====================================================
        S_CAP: begin
          // �Է� �ȼ��� in_valid �޽� ���� 1���� ���´�.
          if (in_valid) begin
            fb[wr_addr] <= in_pixel;
            wr_addr     <= wr_addr + {{(A_W-1){1'b0}},1'b1};
          end

          // ������ �� �Ǵ�: ������ ���� ������ �ȼ����� in_line_last�� 1clk
          // (TB/�������� mp_frame_last�� �ִٸ� �װ��� Ȱ���ص� ��)
          if (ill_rise && (wr_addr == DEPTH-1)) begin
            // ĸó �Ϸ� �� TOP PAD�� ���� (������ �����Ǿ� �־�� ��)
            st         <= S_TOP;
            rd_addr    <= {A_W{1'b0}};
            px_in_line <= 10'd0;
            lines_done <= 7'd0;
          end
        end

        // ====================================================
        // 2) TOP PADDING (PAD lines)
        // ====================================================
        S_TOP: begin
          if (slot_tick) begin
            out_valid  <= 1'b1;
            out_is_pad <= 1'b1;
            out_pixel  <= 8'd0;

            if (px_in_line == W-1) begin
              out_line_last <= 1'b1;
              px_in_line    <= 10'd0;
              if (lines_done == PAD-1) begin
                st         <= S_PAY;
                lines_done <= 7'd0;
              end else begin
                lines_done <= lines_done + 7'd1;
              end
            end else begin
              px_in_line <= px_in_line + 10'd1;
            end
          end
        end

        // ====================================================
        // 3) PAYLOAD REPLAY (HIN lines)
        // ====================================================
        S_PAY: begin
          if (slot_tick) begin
            out_valid  <= 1'b1;
            out_is_pad <= 1'b0;
            out_pixel  <= fb[rd_addr];
            rd_addr    <= rd_addr + {{(A_W-1){1'b0}},1'b1};

            if (px_in_line == W-1) begin
              out_line_last <= 1'b1;
              px_in_line    <= 10'd0;
              if (lines_done == HIN-1) begin
                st         <= S_BOT;
                lines_done <= 7'd0;
              end else begin
                lines_done <= lines_done + 7'd1;
              end
            end else begin
              px_in_line <= px_in_line + 10'd1;
            end
          end
        end

        // ====================================================
        // 4) BOTTOM PADDING (PAD lines)
        // ====================================================
        S_BOT: begin
          if (slot_tick) begin
            out_valid  <= 1'b1;
            out_is_pad <= 1'b1;
            out_pixel  <= 8'd0;

            if (px_in_line == W-1) begin
              out_line_last <= 1'b1;
              px_in_line    <= 10'd0;
              if (lines_done == PAD-1) begin
                out_frame_last <= 1'b1;   // �������� ������ �ȼ�
                // ���� ������ �غ� (�ٽ� CAP����)
                st         <= S_CAP;
                wr_addr    <= {A_W{1'b0}};
                rd_addr    <= {A_W{1'b0}};
                lines_done <= 7'd0;
              end else begin
                lines_done <= lines_done + 7'd1;
              end
            end else begin
              px_in_line <= px_in_line + 10'd1;
            end
          end
        end

        default: st <= S_CAP;
      endcase
    end
  end

endmodule


