// quantize_s8.v  (ZERO_POINT ���� ����ȭ, PAD=0 ����)
module quantize_s8 #(
  parameter signed [7:0] ZERO_POINT = 8'sd128
)(
  input  wire             clk,
  input  wire             srst,            // active-HIGH
  // in (valid-gated stream)
  input  wire             in_valid,
  input  wire      [7:0]  in_pixel,        // u8
  input  wire             in_line_last,
  input  wire             in_frame_last,
  input  wire             in_is_pad,       // 1 = pad �ȼ�

  // out
  output reg              out_valid,
  output reg signed [7:0] out_pixel,       // s8
  output reg              out_line_last,
  output reg              out_frame_last,
  output reg              out_is_pad
);

  // ������ 1�� (valid�� �Բ� ����)
  reg             vld_ff;
  reg      [7:0]  pix_ff;
  reg             ll_ff, fl_ff;
  reg             pad_ff;

  always @(posedge clk) begin
    if (srst) begin
      vld_ff <= 1'b0;
      pix_ff <= 8'd0;
      ll_ff  <= 1'b0;
      fl_ff  <= 1'b0;
      pad_ff <= 1'b0;
    end else begin
      vld_ff <= in_valid;
      if (in_valid) begin
        pix_ff <= in_pixel;
        ll_ff  <= in_line_last;
        fl_ff  <= in_frame_last;
        pad_ff <= in_is_pad;          // �� PAD �÷��׸� valid�� �Բ� ���ø�
      end else begin
        // valid�� 0�� �� '���� �� ����'(���� ä���)
        ll_ff  <= 1'b0;
        fl_ff  <= 1'b0;
        pad_ff <= 1'b0;
      end
    end
  end

  // ������ 2��: ���� ����ȭ + PAD=0 ����
  always @(posedge clk) begin
    if (srst) begin
      out_valid      <= 1'b0;
      out_pixel      <= 8'sd0;
      out_line_last  <= 1'b0;
      out_frame_last <= 1'b0;
      out_is_pad     <= 1'b0;
    end else begin
      out_valid      <= vld_ff;
      out_line_last  <= vld_ff ? ll_ff  : 1'b0;  // �� valid�� ����Ʈ
      out_frame_last <= vld_ff ? fl_ff  : 1'b0;  // �� valid�� ����Ʈ
      out_is_pad     <= vld_ff ? pad_ff : 1'b0;  // �� PAD �÷��� ����

      if (vld_ff) begin
        // �� PAD�� ������ 0. �׷��� ������ (u8 - ZERO_POINT)
        if (pad_ff) begin
          out_pixel <= 8'sd0;
        end else begin
          // u8 -> s9�� Ȯ�� �� ZERO_POINT ���� (wrap ������)
          out_pixel <= $signed({1'b0, pix_ff}) - $signed(ZERO_POINT);
        end
      end
    end
  end
endmodule
